
module anemoVER_1_0 (
	clk_clk,
	in_freq_anemometre_beginbursttransfer,
	reset_reset_n,
	test_export);	

	input		clk_clk;
	input		in_freq_anemometre_beginbursttransfer;
	input		reset_reset_n;
	output	[7:0]	test_export;
endmodule
